Baker Chapter 6 Figure 6.11 - NMOS Curve Trace 

* FET model using built-in default parameters for BSIM4
.model nm1 nmos level=54 version=4.8.1
.model pm1 pmos level=54 version=4.8.1

* 
* IMPORTANT: We are running with this line in the .spiceinit file:
* 
* optran 0 0 0 100p 50n 0 ; Don't use DC operating point, but transient op
*

Vds vds 0 dc 2
Vgs vgs 0 dc 3

* NMOS (drain, gate, source, body).
M1 vds vgs 0 0 nm1 W=10 L=1

.control
destroy all
.options savecurrents
.option scale=1u 
dc vds 0 3 0.5 vgs 0 2 0.5
plot -1*i(vds)
.endc
.end
