NMOS Demo #1 using Skywater 130 model

.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

Vdd vdd 0 1.8
Vss vss 0 0
* Fixed Vgs
Vgs in 0 1.8

* Notice that the MOSFET is represented here as a subcircuit (starts with X!)
* NMOS pin convention: drain, gate, source, body.
XMn1 vdd in vss vss sky130_fd_pr__nfet_01v8_lvt 
+ L=0.15 W=1 nf=1 
+ sa=0 sb=0 sd=0 mult=1 m=1
+ ad='int((nf+1)/2) * W/nf * 0.29' 
+ as='int((nf+2)/2) * W/nf * 0.29' 
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' 
+ nrd='0.29 / W' 
+ nrs='0.29 / W' 

.control
* Transient analysis
tran 100p 1000n 10n
set xbrushwidth=2
plot -1 * i(vdd)
.endc
.end
