voltage divider
V1 in 0 dc 0 PULSE (0 1 1u 1u 1u 1 1)
*V1 in 0 1
R1 in out 1k
R2 out 0 2k
.end


