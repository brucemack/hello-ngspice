inverter example circuit for control language tutorial
* file inv-example2.cir

* the power supply 
Vcc cc 0 1

* the input signal for dc and tran simulation
Vin in 0 dc 0 pulse (0 1 95n 2n 2n 90n 180n)

* the circuit
Mn1 out in 0 0 nm W=2u L=0.18u
Mp1 out in cc cc pm W=4u L=0.18u

* model and model parameters (we use the built-in default parameters for BSIM4)
.model nm nmos level=14 version=4.8.1
.model pm pmos level=14 version=4.8.1

* control language script
.control
tran 100p 500n               ; simulation command 1
set xbrushwidth=2
plot v(in) v(out)
write $inputdir/outtran.out v(in) v(out)
reset
dc vin 0 1 0.01              ; simulation command 2
plot v(out)                  ; v(in) not required because it is the x axis already
write $inputdir/outdc.out v(out)
.endc
.end
